library IEEE;
use IEEE.std_logic_1164.all;

entity i_cache is
port( 	in_add : in std_logic_vector(4 downto 0);
	output: out std_logic_vector(31 downto 0)
	);

end i_cache;

architecture behav of i_cache is
begin
	process(in_add)
	begin
		case in_add is
	when "00001" =>
		output <= "00000000000000000000000000000000";
	when "00010" =>
		output <= "00000000000000000000000000000000";
	when "00011" =>
		output <= "00000000000000000000000000000000";
	when "00100" =>
		output <= "00000000000000000000000000000000";
	when "00101" =>
		output <= "00000000000000000000000000000000";
	when "00110" =>
		output <= "00000000000000000000000000000000";
	when "00111" =>
		output <= "00000000000000000000000000000000";
	when "01000" =>
		output <= "00000000000000000000000000000000";
	when "01001" =>
		output <= "00000000000000000000000000000000";
	when "01010" =>
		output <= "00000000000000000000000000000000";
	when "01011" =>
		output <= "00000000000000000000000000000000";
	when "01100" =>
		output <= "00000000000000000000000000000000";
	when "01101" =>
		output <= "00000000000000000000000000000000";
	when "01110" =>
		output <= "00000000000000000000000000000000";
	when "01111" =>
		output <= "00000000000000000000000000000000";
	when "10000" =>
		output <= "00000000000000000000000000000000";
	when "10001" =>
		output <= "00000000000000000000000000000000";
	when "10010" =>
		output <= "00000000000000000000000000000000";
	when "10011" =>
		output <= "00000000000000000000000000000000";
	when "10100" =>
		output <= "00000000000000000000000000000000";
	when "10101" =>
		output <= "00000000000000000000000000000000";
	when "10110" =>
		output <= "00000000000000000000000000000000";
	when "10111" =>
		output <= "00000000000000000000000000000000";
	when "11000" =>
		output <= "00000000000000000000000000000000";
	when "11001" =>
		output <= "00000000000000000000000000000000";
	when "11010" =>
		output <= "00000000000000000000000000000000";
	when "11011" =>
		output <= "00000000000000000000000000000000";
	when "11100" =>
		output <= "00000000000000000000000000000000";
	when "11101" =>
		output <= "00000000000000000000000000000000";
	when "11110" =>
		output <= "00000000000000000000000000000000";
	when others =>
		output <= "00000000000000000000000000000000";
		end case;	
	end process;
end behav;
